
",{gut*
"r$